* NMOS with pull up resistor

V01 1 0 0.8V
V02 2 0 5V

R23 2 3 R=1000

M310 3 1 0 0 t_model

.OP

.END
