* Simple RC circuit

V01 1 0 EXP( 0.0 3.0 0.0 2n 10n 4n)

R12 1 2 R=1000
C20 2 0 C=1p

.TRAN 40n 1n

.END
