* Simple RL circuit

V01 1 0 3V

R12 1 2 R=1000
L20 2 0 L=1n

*.OP
.TRAN 40m 1m

.END
