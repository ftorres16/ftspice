*Basic test

V1 1 0 4000mV

R12 1 2 R=2200
R20 2 0 R=2.2k

.END
