* Simple RL circuit

V01 1 0 3A

R12 1 2 R=1000
L20 2 0 L=1

.OP
.TRAN 0 1 1m

.END
