* Basic test - Current Divider

I1 1 0 10mA

R10a 1 0 R=2200
R10b 1 0 R=2.2k

.END
