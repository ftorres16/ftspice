*Proj 1

V50 5 0 2V
V76 7 6 2V
V32 3 2 0.2V

I1 6 0 1mA
I2 8 4 1mA

R1 5 1 R=1.5
R2 5 2 R=50
R3 5 6 R=0.1
R4 1 2 R=1
R5 2 6 R=1.5
R6 3 4 R=0.1
R7 4 0 R=10
R8 8 0 R=1000

.OP

.END
