* Basic test - R-D
V1 1 0 4000mV

R12 1 2 R=2200
D20 0 2 d_model

.END
