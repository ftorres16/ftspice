* NPN with pull up resistor

V01 1 0 0.8V
V02 2 0 3V

R23 2 3 R=640
R14 1 4 R=10

Q310 3 4 0 0 q_model

.OP

.END
