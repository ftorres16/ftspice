* Simple RC circuit

I01 1 0 SIN( 0.0 3.0m 100M )

R10 1 0 R=100
C10 1 0 C=10p

.TRAN 0 40n 1n

.END
